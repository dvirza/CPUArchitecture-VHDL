LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package aux_package is
-----------------------------------------------------------------
	component top is
		generic (
			n : integer := 8 );
		port(
			rst,ena,clk : in std_logic
			
		);
	end component;
-----------------------------------------------------------------
	component Adder IS
		GENERIC (n : integer := 16);
		PORT ( a, b: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
		       cin: IN STD_LOGIC;
               s: OUT STD_LOGIC_VECTOR (n-1 DOWNTO 0);
		       cout: OUT STD_LOGIC);
	END component;
-----------------------------------------------------------------
	component aluCore is
			GENERIC (
				n: integer:=8;
				Dwidth: integer:=16;
				opwidth: integer:=4
				);
			port(	srcA,srcB: 	 	   in std_logic_vector(Dwidth-1 downto 0);
				opc: 		 	   in std_logic_vector(opwidth-1 downto 0);
				aluOut:	     	   out std_logic_vector(Dwidth-1 downto 0);
				cFlag,nFlag,zFlag: out std_logic
			);

	end component;
-----------------------------------------------------------------
	component aluTop is
		GENERIC (
			n: integer:=8;
			Dwidth: integer:=16;
			opwidth: integer:=4
			);
		port(	reg_srcA,wire_srcB: 	 			in std_logic_vector(Dwidth-1 downto 0);
			opc_wire: in std_logic_vector (opwidth-1 downto 0);
			clk, rst, regAin, regCin: in std_logic;
			reg_cOut: 							out std_logic_vector(Dwidth-1 downto 0);
			wire_cFlag, wire_zFlag, wire_nFlag: out std_logic
		);
	end component;
-----------------------------------------------------------------
	component pcWork is
		generic( Dwidth: integer:=16;
		Awidth: integer:=6;
		dept:   integer:=64);
		port(	clk,rst,PCin: 		in std_logic;	
			PCsel : 			in std_logic_vector(1 downto 0);
			IRinReg: 			in std_logic_vector(7 downto 0);
			PCdata: 			out std_logic_vector(Awidth-1 downto 0)
		);
	end component; 
-----------------------------------------------------------------
	component ProgMem is
	generic( Dwidth: integer:=16;
			 Awidth: integer:=6;
			 dept:   integer:=64);
	port(	clk,memEn: in std_logic;	
			WmemData:	in std_logic_vector(Dwidth-1 downto 0);
			WmemAddr,RmemAddr:	
						in std_logic_vector(Awidth-1 downto 0);
			RmemData: 	out std_logic_vector(Dwidth-1 downto 0)
	);
	end component;
-----------------------------------------------------------------
	component dataMem is
		generic( Dwidth: integer:=16;
				Awidth: integer:=6;
				dept:   integer:=64);
		port(	clk,memEn: in std_logic;	
				WmemData:	in std_logic_vector(Dwidth-1 downto 0);
				WmemAddr,RmemAddr:	
							in std_logic_vector(Awidth-1 downto 0);
				RmemData: 	out std_logic_vector(Dwidth-1 downto 0)
		);
	end component;
-----------------------------------------------------------------
	component mod_ProgMem is
		generic( Dwidth: integer:=16;
				Awidth: integer:=6;
				dept:   integer:=64);
		port(	clk, rst, tbWren, pcin, tbActive:        in std_logic;
				pcsel : in std_logic_vector(1 downto 0);
				irinreg : in std_logic_vector(7 downto 0);
				tbAddrIn : in std_logic_vector(Awidth-1 downto 0);
				tbDataIn : in std_logic_vector (Dwidth-1 downto 0);
				dataOut: 	out std_logic_vector(Dwidth-1 downto 0)
		);
	end component;
-----------------------------------------------------------------
	component RF is
		generic( Dwidth: integer:=16;
				opwidth: integer:=4);
		port(	clk,rst,WregEn: in std_logic;	
				WregData:	in std_logic_vector(Dwidth-1 downto 0);
				WregAddr,RregAddr:	
							in std_logic_vector(opwidth-1 downto 0);
				RregData: 	out std_logic_vector(Dwidth-1 downto 0)
		);
		end component;
-----------------------------------------------------------------
end package aux_package;